---------------------------------------------------------------------------------
-- Univ. of Chicago  
--    
--
-- PROJECT:      ANNIE - ACDC
-- FILE:         trigger.vhd
-- AUTHOR:       D. Greenshields
-- DATE:         Sep 2020
--
-- DESCRIPTION:  trigger processes
---------------------------------------------------------------------------------

	
library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use work.defs.all;
use work.components.pulseSync;



entity trigger is
	port(
			clock						: in	clock_type;
			reset						: in	std_logic;   
			systemTime				: in  std_logic_vector(63 downto 0);
			testMode					: in  testMode_type;
			trigSetup				: in	trigSetup_type;
			trigInfo					: out	trigInfo_type;
			acc_trig					: in	std_logic;	-- trig from central card (LVDS)
			sma_trig					: in	std_logic;	-- on-board SMA input
			self_trig				: in	std_logic;	
			sma_validate			: in	std_logic;	-- on-board SMA input
			digitize_request		: out	std_logic;
			transfer_request		: out	std_logic;
			digitize_done			: in	std_logic;
			transfer_enable		: out std_logic;	
			transfer_done			: in	std_logic;
			eventCount				: out	natural;
			timestamp				: out std_logic_vector(63 downto 0);
			validate_pass			: buffer std_logic;
			validate_fail			: buffer std_logic;
			trig_validate			: buffer std_logic;
			validate_clear			: buffer std_logic;
			trig_event				: buffer std_logic;
			trig_clear				: buffer std_logic;
			trig_armed				: out std_logic;	-- used for monitoring/test purposes
			trig_out					: buffer std_logic;
			trig_rate_count		: out natural
			);
end trigger;

architecture vhdl of trigger is





	signal 	sma_trig_z:	std_logic;
	signal 	sma_trig_edge_latch:	std_logic;
	signal 	sma_trig_level_latch:	std_logic;
	signal 	sma_trig_latch:	std_logic;
	signal 	sma_validate_z:	std_logic;
	signal 	sma_validate_latch:	std_logic;
	signal 	sma_validate_edge_latch:	std_logic;
	signal 	sma_validate_level_latch:	std_logic;
	signal 	acc_trig_z:	std_logic;
	signal 	acc_trig_edge_latch:	std_logic;
	signal 	acc_trig_level_latch:	std_logic;
	signal 	acc_trig_latch:	std_logic;
	signal 	acc_validate_z:	std_logic;
	signal 	acc_validate_latch:	std_logic;
	signal 	acc_validate_edge_latch:	std_logic;
	signal 	acc_validate_level_latch:	std_logic;
	signal 	self_trig_z:	std_logic;
	signal 	self_trig_latch:	std_logic;
	signal 	self_trig_edge_latch:	std_logic;
	signal 	self_trig_level_latch:	std_logic;
	signal	self_trig_combined:	std_logic;
	signal	self_trig_sum: natural range 0 to 31;
	signal 	self_trig_enable:	std_logic;
	signal	self_trig_reg: array6;
	signal	self_trig_psec_chip_sum: array6;
	signal 	pps_trig_enable:	std_logic;
	signal	psec_chip_sum: natArray4;
	signal 	selfTrig_rateCount_z: selfTrig_rateCount_array;
	signal	rateCount_valid: std_logic;
	signal	rateCount_valid_z: std_logic;
	signal 	trig_detect:	std_logic;
	signal 	trig_detect_z:	std_logic;
	signal	trig_z2: std_logic;
	signal	trig_detect_arm: std_logic;
	signal	trig_detect_arm_z: std_logic;
	signal	trig_detect_arm_z2: std_logic;
	signal	trig_validate_z:	std_logic;
	signal 	trig_holdoff:	std_logic;
	signal	prev_mode: natural;
	signal	trig_common: std_logic;
	signal	trig_common_z: std_logic;
	signal	resetRequest: std_logic;
	signal	trig_clocked: std_logic;
	signal	trig_clocked_z: std_logic;
	signal	shift_reg: std_logic_vector(7 downto 0);
	signal	trig_sync: std_logic;
	signal	trig_delayed: std_logic;
	signal	sw_trig_enable: std_logic;
	signal	acdc_sma_trig_enable: std_logic;
	signal	acc_sma_trig_enable: std_logic;
	signal	acdc_sma_validate_enable: std_logic;
	signal	acc_sma_validate_enable: std_logic;
	signal	timestamp_z: std_logic_vector(63 downto 0);
	signal	validate_fail_z: std_logic;
	signal	validate_pass_z: std_logic;
	signal	valid_window_end: natural range 0 to 65535;
	
	
	
	
	
begin  



-- brief description:
---------------------
-- A trigger is detected which has different sources depending on the mode:-
--
-- sma input
-- acc via lvds
-- self trigger (generated by psec4 chips when signal level exceeds threshold on a number of channels
--
-- For some modes a validation signal must also be received within a certain time of the trigger
-- This can come from sma input or acc
--









------------------
-- TRIG DETECT
------------------

-- clock the trigger signal and detect a rising edge on it
-- then immediately get a timestamp of when the trigger occurred
-- and generate a flag to initiate subsequent (less time critical) processes
TRIG_DETECTOR: process(clock.x8)
variable t: std_logic;
variable trig_detect_enable: std_logic;
begin
	if (rising_edge(clock.x8)) then		
		
		-- rising edge on 'trig detect arm' enables trigger detection
		-- we only want to detect one trigger at a time and then wait until it has been fully processed
		trig_detect_arm_z <= trig_detect_arm;
		trig_detect_arm_z2 <= trig_detect_arm_z;
		if (trig_detect_arm_z = '1' and trig_detect_arm_z2 = '0') then
			trig_detect_enable := '1';
		end if;
		
		t := '0';
		trig_z2 <= trig_common_z;
		if (trig_detect_enable = '1') then
			if (trig_z2 = '0' and trig_common_z = '1') then		-- rising edge
				t := '1';
				trig_detect_enable := '0';
				timestamp_z <= systemTime;
			end if;
		end if;
		
		trig_detect <= t;
		trig_armed <= trig_detect_enable;
		
	end if;
end process;


-- synchronize trig detect to sys clock
SYNC0: pulseSync port map (clock.x8, clock.sys, trig_detect, trig_detect_z);
	


	
	
	
	
-------------------------
-- VALIDATE CHECK
-------------------------

-- checks if a validation signal was received within the specified time window
VALIDATE_WINDOW_LATCH: process(clock.sys)
variable t: natural range 0 to 65535;
variable busy: boolean;
begin
	if (rising_edge(clock.sys)) then		
		
		trig_validate_z <= trig_validate;
		
		valid_window_end <= trigSetup.valid_window_start + trigSetup.valid_window_len;
		
		if (trig_detect_z = '1') then
		
			validate_clear <= '1';		-- clear the validation latches. These remain in reset until the window start
			validate_fail_z <= '0';
			validate_pass_z <= '0';
			busy := true;
			t := 1;			-- time since the trigger pulse
		
		elsif (busy) then
		
			t := t + 1;
			if (t >= valid_window_end) then
				validate_fail_z <= '1';		-- end of window; no valid signal was received
				busy := false;
			elsif (t >= trigSetup.valid_window_start) then
				validate_clear <= '0';		-- enable the validation latches
				if (trig_validate_z = '1') then	-- a valid signal was received
					validate_pass_z <= '1';
					busy := false;
				end if;
			end if;
			
		end if;				
			
	
	end if;
end process;

	





	

---------------------------------------
-- TRIGGER CONTROL STATE MACHINE
---------------------------------------

TRIG_CTRL: process(clock.sys)
type state_type is (IDLE, VALIDATE, DIGITIZE_BEGIN, DIGITIZE_WAIT, WAIT_FOR_SYSTEM, TRANSFER, TRIG_RESET);
variable state: state_type;
variable transfer_en: boolean;	-- allow transfer of data to acc
variable trig_en : std_logic_vector(4 downto 0);
variable validate_en : std_logic_vector(1 downto 0);
begin
	if (rising_edge(clock.sys)) then
	
		-- synchronize valid check signals to sys clock
		validate_pass <= validate_pass_z;
		validate_fail <= validate_fail_z;
		
		prev_mode <= trigSetup.mode;
		if (prev_mode /= trigSetup.mode) then state := TRIG_RESET; end if;			
		if (trigSetup.resetReq = '1') then state := TRIG_RESET; end if;		-- a trig reset request from acc
				
		
		if (reset = '1' or trigSetup.eventAndTime_reset = '1') then 


			transfer_en := false;
			trig_holdoff <= '0';
			trig_clear <= '1';
			trig_event <= '0';
			
			-- mode control
			sw_trig_enable <= '0'; 
			acdc_sma_trig_enable <= '0';
			acc_sma_trig_enable <= '0';
			self_trig_enable <= '0';
			
			state := TRIG_RESET;
			eventCount <= 0;
		

		else
		

			if (trigSetup.transferEnableReq = '1') then transfer_en := true; end if;
			if (trigSetup.transferDisableReq = '1') then transfer_en := false; end if;

			case state is
			
			
			
				when TRIG_RESET =>
				
					trig_clear <= '1';		-- clear the latches
					trig_holdoff <= '0';		-- enable the trigger sources
					trig_event <= '0';
					trig_detect_arm <= '0';
					state := IDLE;
	
	
	
	
				when IDLE =>		-- waiting for a new trigger signal
				
					
					trig_detect_arm <= '1';		-- enable trigger detection
					trig_clear <= '0';		-- enable the trigger latches


					-- the following switch enables the trigger sources and validation sources
					case trigSetup.mode is
					
						-- trig_en 		:= self & acdc & acc & sw & pps
						-- validate_en	:= acdc & acc						
						when 0 => trig_en := "00000"; validate_en := "00";	-- trigger off
						when 1 => trig_en := "00010"; validate_en := "00";	-- software trigger (from acc)
						when 2 => trig_en := "00100"; validate_en := "00";	-- sma trigger (ACC)
						when 3 => trig_en := "01000"; validate_en := "00";	-- sma trigger (ACDC)
						when 4 => trig_en := "10000"; validate_en := "00";	-- self trigger 
						when 5 => trig_en := "10000"; validate_en := "01";	-- self trigger with sma validation (ACC)
						when 6 => trig_en := "10000"; validate_en := "10";	-- self trigger with sma validation (ACDC)
						when 7 => trig_en := "00100"; validate_en := "10";	-- sma trigger (ACC) with sma validation (ACDC)
						when 8 => trig_en := "01000"; validate_en := "01";	-- sma trigger (ACDC) with sma validation (ACC)
						when 9 => trig_en := "00001"; validate_en := "00";	-- pps trigger (from ACC)
						when others => trig_en := "00000"; validate_en := "00";	-- trigger off

						
					end case;					
					
					pps_trig_enable 			<= trig_en(0);
					sw_trig_enable 			<= trig_en(1); 
					acc_sma_trig_enable 		<= trig_en(2);
					acdc_sma_trig_enable 	<= trig_en(3);
					self_trig_enable 			<= trig_en(4);
					
					acc_sma_validate_enable 	<= validate_en(0);
					acdc_sma_validate_enable 	<= validate_en(1);
					
					if (trig_detect_z = '1') then		-- a trigger rising edge occurred 
			
						timestamp <= timestamp_z;	-- sync the timestamp output to the system clock
						trig_holdoff <= '1';		-- prevent any more triggers while this is high
						
						if (validate_en /= "00") then		-- validation required
							state := VALIDATE;
						elsif (trig_en /= "0000") then	-- no validation required
							state := DIGITIZE_BEGIN;						
						end if;
					
					
					end if;
				
				
				
				
				
				when VALIDATE =>		-- trigger was detected (PSEC4s have captured the data), now wait for validation signals within a specified time window		
					
					if (validate_pass = '1') then 	-- a coincident signal was received, the trig event is valid
						state := DIGITIZE_BEGIN;		
					elsif (validate_fail = '1') then		-- reached the end of the validation window, no valid signal was received - discard the trigger event
						state := TRIG_RESET;			
					end if;					
						
						
								
						
				
				when DIGITIZE_BEGIN =>
				
					eventCount <= eventCount + 1;
					trig_event <= '1';		-- flag used to latch the timestamp and event count externally
					if (testMode.trig_noTransfer = '1') then 
						state := TRIG_RESET;
					else
						digitize_request <= '1';
						state := DIGITIZE_WAIT;
					end if;
				
				
				
				
				when DIGITIZE_WAIT =>
				
					trig_event <= '0';
					digitize_request <= '0';
					if (digitize_done = '1') then 
						state := WAIT_FOR_SYSTEM;		-- don't send data to acc yet as it may be busy processing the previous data
					end if;
						
				
				
				
				when WAIT_FOR_SYSTEM =>		-- wait until the 'transfer enable' signal appears		
					
					if (transfer_en) then			-- transfer enable means one set of data may be transferred
						transfer_request <= '1';
						transfer_en := false;
						state := TRANSFER;
					end if;
				
				
				
				
				when TRANSFER =>		-- transfer data to the acc
				
					transfer_request <= '0';
					if (transfer_done = '1') then		-- data was transferred, now reset ready for the next trigger
						state := TRIG_RESET;
					end if;
					
					
				
				

						
			end case;
				
				
		end if;
		
		if (transfer_en) then transfer_enable <= '1'; else transfer_enable <= '0'; end if;
		
	end if;
	
end process;




	
	
	
	
	
	
	
---------------------------------------
-- ACDC SMA TRIGGER 
---------------------------------------


-- polarity invert option
sma_trig_z <= sma_trig xor trigSetup.sma_invert;		-- 1 = falling edge or low level; 0 = rising edge or high level



-- Edge detect
SMA_TRIG_EDGE_DETECT: process(sma_trig_z, trig_clear, acdc_sma_trig_enable, trig_holdoff)
begin
	if (trig_clear = '1') then
		sma_trig_edge_latch <= '0';
	elsif (rising_edge(sma_trig_z) and acdc_sma_trig_enable = '1' and trig_holdoff = '0') then
		sma_trig_edge_latch <= '1';
	end if;
end process;


-- Level detect
SMA_TRIG_LEVEL_DETECT: process(sma_trig_z, trig_clear, acdc_sma_trig_enable, trig_holdoff)
begin
	if (trig_clear = '1') then
		sma_trig_level_latch <= '0';
	elsif (sma_trig_z = '1' and acdc_sma_trig_enable = '1' and trig_holdoff = '0') then
		sma_trig_level_latch <= '1';
	end if;
end process;
	


-- output select
sma_trig_latch <= sma_trig_edge_latch when (trigSetup.sma_detect_mode = '0') else sma_trig_level_latch;





---------------------------------------
-- ACC TRIGGER 
---------------------------------------
-- trigger coming from acc via lvds
-- This could be from software, from the SMA input on the acc board or from the pps input
-- If from software or pps, use fixed rising-edge-triggered option


-- polarity invert option (only for acc sma option, not acc sw option)
acc_trig_z <= acc_trig xor (trigSetup.acc_invert and acc_sma_trig_enable);		-- 1 = falling edge or low level; 0 = rising edge or high level



-- Edge detect
ACC_TRIG_EDGE_DETECT: process(acc_trig_z, trig_clear, acc_sma_trig_enable, sw_trig_enable, trig_holdoff)
begin
	if (trig_clear = '1') then
		acc_trig_edge_latch <= '0';
	elsif (rising_edge(acc_trig_z) and (acc_sma_trig_enable = '1' or sw_trig_enable = '1' or pps_trig_enable = '1') and trig_holdoff = '0') then
		acc_trig_edge_latch <= '1';
	end if;
end process;


-- Level detect
ACC_TRIG_LEVEL_DETECT: process(acc_trig_z, trig_clear, acc_sma_trig_enable, trig_holdoff)
begin
	if (trig_clear = '1') then
		acc_trig_level_latch <= '0';
	elsif (acc_trig_z = '1' and acc_sma_trig_enable = '1' and trig_holdoff = '0') then
		acc_trig_level_latch <= '1';
	end if;
end process;



-- output select
acc_trig_latch <= acc_trig_level_latch when (trigSetup.acc_detect_mode = '1' and acc_sma_trig_enable = '1')
	else acc_trig_edge_latch;






---------------------------------------
-- SELF TRIGGER 
---------------------------------------



-- Edge detect
SELF_TRIG_EDGE_DETECT: process(self_trig, trig_clear, self_trig_enable, trig_holdoff)
begin
	if (trig_clear = '1') then
		self_trig_edge_latch <= '0';
	elsif (rising_edge(self_trig) and self_trig_enable = '1' and trig_holdoff = '0') then
		self_trig_edge_latch <= '1';
	end if;
end process;


-- Level detect
SELF_TRIG_LEVEL_DETECT: process(self_trig, trig_clear, self_trig_enable, trig_holdoff)
begin
	if (trig_clear = '1') then
		self_trig_level_latch <= '0';
	elsif (self_trig = '1' and self_trig_enable = '1' and trig_holdoff = '0') then
		self_trig_level_latch <= '1';
	end if;
end process;


-- output select
self_trig_latch <= self_trig_edge_latch when (trigSetup.selfTrig_detect_mode = '0') else self_trig_level_latch;





---------------------------------------
-- TRIGGER OUT
---------------------------------------

-- common trigger signal 
trig_common <= (sma_trig_latch or acc_trig_latch or self_trig_latch) and trigSetup.enable;


CLOCKED_TRIG_GEN: process(clock.x8)
begin
	if (rising_edge(clock.x8)) then
		trig_common_z <= trig_common;		-- synchronize to fast clock
	end if;
end process;


TRIG_MULTIPLEXER: process(trigSetup, trig_common_z, trig_common)
begin
	if (trigSetup.use_clocked_trig = '1') then
		trig_out <= trig_common_z;
	else
		trig_out <= trig_common;
	end if;
end process;










---------------------------------------
-- ACDC SMA VALIDATE 
---------------------------------------


-- polarity invert option
sma_validate_z <= sma_validate xor trigSetup.sma_invert;		-- 1 = falling edge or low level; 0 = rising edge or high level



-- Edge detect
SMA_VALIDATE_EDGE_DETECT: process(sma_validate_z, validate_clear, acdc_sma_validate_enable)
begin
	if (validate_clear = '1') then
		sma_validate_edge_latch <= '0';
	elsif (rising_edge(sma_validate_z) and acdc_sma_validate_enable = '1') then
		sma_validate_edge_latch <= '1';
	end if;
end process;


-- Level detect
SMA_VALIDATE_LEVEL_DETECT: process(sma_validate_z, validate_clear, acdc_sma_validate_enable)
begin
	if (validate_clear = '1') then
		sma_validate_level_latch <= '0';
	elsif (sma_validate_z = '1' and acdc_sma_validate_enable = '1') then
		sma_validate_level_latch <= '1';
	end if;
end process;


-- output select
sma_validate_latch <= sma_validate_edge_latch when (trigSetup.sma_detect_mode = '0') else sma_validate_level_latch;





---------------------------------------
-- ACC SMA VALIDATE 
---------------------------------------
-- validation coming from the SMA connector on the acc board via lvds


-- polarity invert option
acc_validate_z <= acc_trig xor trigSetup.acc_invert;		-- 1 = falling edge or low level; 0 = rising edge or high level



-- Edge detect
ACC_VALIDATE_EDGE_DETECT: process(acc_validate_z, validate_clear, acc_sma_validate_enable)
begin
	if (validate_clear = '1') then
		acc_validate_edge_latch <= '0';
	elsif (rising_edge(acc_validate_z) and acc_sma_validate_enable = '1') then
		acc_validate_edge_latch <= '1';
	end if;
end process;


-- Level detect
ACC_VALIDATE_LEVEL_DETECT: process(acc_validate_z, validate_clear, acc_sma_validate_enable)
begin
	if (validate_clear = '1') then
		acc_validate_level_latch <= '0';
	elsif (acc_validate_z = '1' and acc_sma_validate_enable = '1') then
		acc_validate_level_latch <= '1';
	end if;
end process;



-- output select
acc_validate_latch <= acc_validate_edge_latch when (trigSetup.acc_detect_mode = '0') else acc_validate_level_latch;






---------------------------------------
-- TRIGGER VALIDATE
---------------------------------------

-- common trigger validation signal
trig_validate <= sma_validate_latch or acc_validate_latch;












------------------
-- TRIG INFO
------------------
-- read back as part of the psec data frame
-- serves as confirmation of the trigger setup status

--
trigInfo(0,0) <= x"EEEE";
trigInfo(0,1)(3 downto 0) <= std_logic_vector(to_unsigned(trigSetup.mode, 4));
trigInfo(0,1)(15 downto 4) <= std_logic_vector(to_unsigned(trigSetup.valid_window_start, 12));

trigInfo(0,2) <= x"0" & std_logic_vector(to_unsigned(trigSetup.valid_window_len, 12));

trigInfo(0,3)(1 downto 0) <= trigSetup.sma_invert & trigSetup.sma_detect_mode;
trigInfo(0,3)(3 downto 2) <= trigSetup.acc_invert & trigSetup.acc_detect_mode;
trigInfo(0,3)(5 downto 4) <= trigSetup.selfTrig_sign & trigSetup.selfTrig_detect_mode;
trigInfo(0,3)(15 downto 6) <= "00000" & std_logic_vector(to_unsigned(trigSetup.selfTrig_coincidence_min, 5));
trigInfo(0,4) <= x"EEEE";

--
trigInfo(1,0) <= "0000000000" & trigSetup.selfTrig_mask(0);
trigInfo(1,1) <= "0000000000" & trigSetup.selfTrig_mask(1);
trigInfo(1,2) <= "0000000000" & trigSetup.selfTrig_mask(2);
trigInfo(1,3) <= "0000000000" & trigSetup.selfTrig_mask(3);
trigInfo(1,4) <= "0000000000" & trigSetup.selfTrig_mask(4);

--
trigInfo(2,0) <= x"0" & std_logic_vector(to_unsigned(trigSetup.selfTrig_threshold(0), 12));
trigInfo(2,1) <= x"0" & std_logic_vector(to_unsigned(trigSetup.selfTrig_threshold(1), 12));
trigInfo(2,2) <= x"0" & std_logic_vector(to_unsigned(trigSetup.selfTrig_threshold(2), 12));
trigInfo(2,3) <= x"0" & std_logic_vector(to_unsigned(trigSetup.selfTrig_threshold(3), 12));
trigInfo(2,4) <= x"0" & std_logic_vector(to_unsigned(trigSetup.selfTrig_threshold(4), 12));








------------------------------
-- TRIGGER RATE COUNTER
------------------------------
-- count the number of trig events in one second 

RATE_COUNT_GEN: process(clock.sys)
variable count: natural;
variable t: natural;
begin
	if (rising_edge(clock.sys)) then
		
		if (reset = '1' or trigSetup.eventAndTime_reset = '1') then
		
			t := 0;
			count := 0;
			trig_rate_count <= 0;
			
			
		else
		
		
			if (trig_event = '1') then
				if (count < trigRate_MaxCount) then count := count + 1; end if;
			end if;				
			
			t := t + 1;		-- clock cycle counter
			 
			if (t = 40000000) then		-- after 1 second record the count and then reset 

				t := 0;
				trig_rate_count <= count;
				count := 0;
				
			end if;
			
		end if;
		
	end if;
end process;






	
end vhdl;






