
module clockSwitch (
	inclk1x,
	inclk0x,
	clkselect,
	outclk);	

	input		inclk1x;
	input		inclk0x;
	input		clkselect;
	output		outclk;
endmodule
